
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.array_generate.all;

entity blocks is
	port(
		clk          : in std_logic;
		LvL_sel : in std_logic_vector(1 downto 0);
		game_state   : in state;
		block_dimensions   : out block_array);
end blocks;

architecture Behavioral of blocks is
begin
    --- In this process, the blocks are assigned to their individual pixel positions ---
    --- As there are 4 levels, in each level there is a different design of the blocks ---
	LvL_Blocks: process(clk, game_state)
	begin
		if rising_edge(clk) and game_state = waiting then
			case LvL_sel is
				when "00" =>
					block_dimensions(0)(0) <= 240;  block_dimensions(16)(0) <= 220;
					block_dimensions(0)(1) <= 0;    block_dimensions(16)(1) <= 0;  
					block_dimensions(0)(2) <= 260;  block_dimensions(16)(2) <= 240;
					block_dimensions(0)(3) <= 40;   block_dimensions(16)(3) <= 40; 
					block_dimensions(1)(0) <= 240;  block_dimensions(17)(0) <= 220;
					block_dimensions(1)(1) <= 40;   block_dimensions(17)(1) <= 40; 
					block_dimensions(1)(2) <= 260;  block_dimensions(17)(2) <= 240;
					block_dimensions(1)(3) <= 80;   block_dimensions(17)(3) <= 80; 
					block_dimensions(2)(0) <= 240;  block_dimensions(18)(0) <= 220;
					block_dimensions(2)(1) <= 80;   block_dimensions(18)(1) <= 80; 
					block_dimensions(2)(2) <= 260;  block_dimensions(18)(2) <= 240;
					block_dimensions(2)(3) <= 120;  block_dimensions(18)(3) <= 120;
					block_dimensions(3)(0) <= 240;  block_dimensions(19)(0) <= 220;
					block_dimensions(3)(1) <= 120;  block_dimensions(19)(1) <= 120;
					block_dimensions(3)(2) <= 260;  block_dimensions(19)(2) <= 240;
					block_dimensions(3)(3) <= 160;  block_dimensions(19)(3) <= 160;
					block_dimensions(4)(0) <= 240;  block_dimensions(20)(0) <= 220;
					block_dimensions(4)(1) <= 160;  block_dimensions(20)(1) <= 160;
					block_dimensions(4)(2) <= 260;  block_dimensions(20)(2) <= 240;
					block_dimensions(4)(3) <= 200;  block_dimensions(20)(3) <= 200;
					block_dimensions(5)(0) <= 240;  block_dimensions(21)(0) <= 220;
					block_dimensions(5)(1) <= 200;  block_dimensions(21)(1) <= 200;
					block_dimensions(5)(2) <= 260;  block_dimensions(21)(2) <= 240;
					block_dimensions(5)(3) <= 240;  block_dimensions(21)(3) <= 240;
					block_dimensions(6)(0) <= 240;  block_dimensions(22)(0) <= 220;
					block_dimensions(6)(1) <= 240;  block_dimensions(22)(1) <= 240;
					block_dimensions(6)(2) <= 260;  block_dimensions(22)(2) <= 240;
					block_dimensions(6)(3) <= 280;  block_dimensions(22)(3) <= 280;
					block_dimensions(7)(0) <= 240;  block_dimensions(23)(0) <= 220;
					block_dimensions(7)(1) <= 280;  block_dimensions(23)(1) <= 280;
					block_dimensions(7)(2) <= 260;  block_dimensions(23)(2) <= 240;
					block_dimensions(7)(3) <= 320;  block_dimensions(23)(3) <= 320;
					block_dimensions(8)(0) <= 240;  block_dimensions(24)(0) <= 220;
					block_dimensions(8)(1) <= 320;  block_dimensions(24)(1) <= 320;
					block_dimensions(8)(2) <= 260;  block_dimensions(24)(2) <= 240;
					block_dimensions(8)(3) <= 360;  block_dimensions(24)(3) <= 360;
					block_dimensions(9)(0) <= 240;  block_dimensions(25)(0) <= 220;
					block_dimensions(9)(1) <= 360;  block_dimensions(25)(1) <= 360;
					block_dimensions(9)(2) <= 260;  block_dimensions(25)(2) <= 240;
					block_dimensions(9)(3) <= 400;  block_dimensions(25)(3) <= 400;
					block_dimensions(10)(0) <= 240; block_dimensions(26)(0) <= 220;
                    block_dimensions(10)(1) <= 400; block_dimensions(26)(1) <= 400;                                            
                    block_dimensions(10)(2) <= 260; block_dimensions(26)(2) <= 240;                                            
                    block_dimensions(10)(3) <= 440; block_dimensions(26)(3) <= 440;                                            
                    block_dimensions(11)(0) <= 240; block_dimensions(27)(0) <= 220;                                            
                    block_dimensions(11)(1) <= 440; block_dimensions(27)(1) <= 440;                                            
                    block_dimensions(11)(2) <= 260; block_dimensions(27)(2) <= 240;                                            
                    block_dimensions(11)(3) <= 480; block_dimensions(27)(3) <= 480;                                            
                    block_dimensions(12)(0) <= 240; block_dimensions(28)(0) <= 220;                                            
                    block_dimensions(12)(1) <= 480; block_dimensions(28)(1) <= 480;                                            
                    block_dimensions(12)(2) <= 260; block_dimensions(28)(2) <= 240;                                            
                    block_dimensions(12)(3) <= 520; block_dimensions(28)(3) <= 520;                                            
                    block_dimensions(13)(0) <= 240; block_dimensions(29)(0) <= 220;                                            
                    block_dimensions(13)(1) <= 520; block_dimensions(29)(1) <= 520;                                            
                    block_dimensions(13)(2) <= 260; block_dimensions(29)(2) <= 240;                                            
                    block_dimensions(13)(3) <= 560; block_dimensions(29)(3) <= 560;                                            
                    block_dimensions(14)(0) <= 240; block_dimensions(30)(0) <= 220;                                            
                    block_dimensions(14)(1) <= 560; block_dimensions(30)(1) <= 560;                                            
                    block_dimensions(14)(2) <= 260; block_dimensions(30)(2) <= 240;                                            
                    block_dimensions(14)(3) <= 600; block_dimensions(30)(3) <= 600;                                            
                    block_dimensions(15)(0) <= 240; block_dimensions(31)(0) <= 220;                                            
                    block_dimensions(15)(1) <= 600; block_dimensions(31)(1) <= 600;                                            
                    block_dimensions(15)(2) <= 260; block_dimensions(31)(2) <= 240;                                            
                    block_dimensions(15)(3) <= 640; block_dimensions(31)(3) <= 640;                                            
                                                                        
                    when "01" =>
					block_dimensions(0)(0) <= 300;  block_dimensions(16)(0) <= 240;
					block_dimensions(0)(1) <= 120;  block_dimensions(16)(1) <= 360;
					block_dimensions(0)(2) <= 320;  block_dimensions(16)(2) <= 260;
					block_dimensions(0)(3) <= 160;  block_dimensions(16)(3) <= 400;
					block_dimensions(1)(0) <= 300;  block_dimensions(17)(0) <= 240;
					block_dimensions(1)(1) <= 360;  block_dimensions(17)(1) <= 480;
					block_dimensions(1)(2) <= 320;  block_dimensions(17)(2) <= 260;
					block_dimensions(1)(3) <= 400;  block_dimensions(17)(3) <= 520;
					block_dimensions(2)(0) <= 300;  block_dimensions(18)(0) <= 240;
					block_dimensions(2)(1) <= 600;  block_dimensions(18)(1) <= 600;
					block_dimensions(2)(2) <= 320;  block_dimensions(18)(2) <= 260;
					block_dimensions(2)(3) <= 640;  block_dimensions(18)(3) <= 640;
					block_dimensions(3)(0) <= 280;  block_dimensions(19)(0) <= 220;
					block_dimensions(3)(1) <= 80;   block_dimensions(19)(1) <= 40; 
					block_dimensions(3)(2) <= 300;  block_dimensions(19)(2) <= 240;
					block_dimensions(3)(3) <= 120;  block_dimensions(19)(3) <= 80; 
					block_dimensions(4)(0) <= 280;  block_dimensions(20)(0) <= 220;
					block_dimensions(4)(1) <= 160;  block_dimensions(20)(1) <= 200;
					block_dimensions(4)(2) <= 300;  block_dimensions(20)(2) <= 240;
					block_dimensions(4)(3) <= 200;  block_dimensions(20)(3) <= 240;
					block_dimensions(5)(0) <= 280;  block_dimensions(21)(0) <= 220;
					block_dimensions(5)(1) <= 320;  block_dimensions(21)(1) <= 280;
					block_dimensions(5)(2) <= 300;  block_dimensions(21)(2) <= 240;
					block_dimensions(5)(3) <= 340;  block_dimensions(21)(3) <= 320;
					block_dimensions(6)(0) <= 280;  block_dimensions(22)(0) <= 220;
					block_dimensions(6)(1) <= 400;  block_dimensions(22)(1) <= 440;
					block_dimensions(6)(2) <= 300;  block_dimensions(22)(2) <= 240;
					block_dimensions(6)(3) <= 440;  block_dimensions(22)(3) <= 480;
					block_dimensions(7)(0) <= 280;  block_dimensions(23)(0) <= 220;
					block_dimensions(7)(1) <= 560;  block_dimensions(23)(1) <= 520;
					block_dimensions(7)(2) <= 300;  block_dimensions(23)(2) <= 240;
					block_dimensions(7)(3) <= 600;  block_dimensions(23)(3) <= 560;
					block_dimensions(8)(0) <= 260;  block_dimensions(24)(0) <= 200;
					block_dimensions(8)(1) <= 40;   block_dimensions(24)(1) <= 80; 
					block_dimensions(8)(2) <= 280;  block_dimensions(24)(2) <= 220;
					block_dimensions(8)(3) <= 80;   block_dimensions(24)(3) <= 120;
					block_dimensions(9)(0) <= 260;  block_dimensions(25)(0) <= 200;
					block_dimensions(9)(1) <= 200;  block_dimensions(25)(1) <= 160;
					block_dimensions(9)(2) <= 280;  block_dimensions(25)(2) <= 220;
					block_dimensions(9)(3) <= 240;  block_dimensions(25)(3) <= 200;
					block_dimensions(10)(0) <= 260; block_dimensions(26)(0) <= 200;
                    block_dimensions(10)(1) <= 280; block_dimensions(26)(1) <= 320;                                            
                    block_dimensions(10)(2) <= 280; block_dimensions(26)(2) <= 220;                                            
                    block_dimensions(10)(3) <= 320; block_dimensions(26)(3) <= 360;                                            
                    block_dimensions(11)(0) <= 260; block_dimensions(27)(0) <= 200;                                            
                    block_dimensions(11)(1) <= 440; block_dimensions(27)(1) <= 400;                                            
                    block_dimensions(11)(2) <= 280; block_dimensions(27)(2) <= 220;                                            
                    block_dimensions(11)(3) <= 480; block_dimensions(27)(3) <= 440;                                            
                    block_dimensions(12)(0) <= 260; block_dimensions(28)(0) <= 200;                                            
                    block_dimensions(12)(1) <= 520; block_dimensions(28)(1) <= 560;                                            
                    block_dimensions(12)(2) <= 280; block_dimensions(28)(2) <= 220;                                            
                    block_dimensions(12)(3) <= 560; block_dimensions(28)(3) <= 600;                                            
                    block_dimensions(13)(0) <= 240; block_dimensions(29)(0) <= 180;                                            
                    block_dimensions(13)(1) <= 0;   block_dimensions(29)(1) <= 160;                                          
                    block_dimensions(13)(2) <= 260; block_dimensions(29)(2) <= 200;                                            
                    block_dimensions(13)(3) <= 40;  block_dimensions(29)(3) <= 200;                                           
                    block_dimensions(14)(0) <= 240; block_dimensions(30)(0) <= 180;                                            
                    block_dimensions(14)(1) <= 120; block_dimensions(30)(1) <= 360;                                            
                    block_dimensions(14)(2) <= 260; block_dimensions(30)(2) <= 200;                                            
                    block_dimensions(14)(3) <= 160; block_dimensions(30)(3) <= 400;                                            
                    block_dimensions(15)(0) <= 240; block_dimensions(31)(0) <= 180;                                            
                    block_dimensions(15)(1) <= 240; block_dimensions(31)(1) <= 600;                                            
                    block_dimensions(15)(2) <= 260; block_dimensions(31)(2) <= 200;                                            
                    block_dimensions(15)(3) <= 280; block_dimensions(31)(3) <= 640;                                            
                                   
                    when "10" =>
					block_dimensions(0)(0) <= 260;  block_dimensions(16)(0) <= 220;
					block_dimensions(0)(1) <= 0;    block_dimensions(16)(1) <= 0;  
					block_dimensions(0)(2) <= 280;  block_dimensions(16)(2) <= 240;
					block_dimensions(0)(3) <= 40;   block_dimensions(16)(3) <= 40; 
					block_dimensions(1)(0) <= 260;  block_dimensions(17)(0) <= 220;
					block_dimensions(1)(1) <= 80;   block_dimensions(17)(1) <= 80; 
					block_dimensions(1)(2) <= 280;  block_dimensions(17)(2) <= 240;
					block_dimensions(1)(3) <= 120;  block_dimensions(17)(3) <= 120;
					block_dimensions(2)(0) <= 260;  block_dimensions(18)(0) <= 220;
					block_dimensions(2)(1) <= 160;  block_dimensions(18)(1) <= 160;
					block_dimensions(2)(2) <= 280;  block_dimensions(18)(2) <= 240;
					block_dimensions(2)(3) <= 200;  block_dimensions(18)(3) <= 200;
					block_dimensions(3)(0) <= 260;  block_dimensions(19)(0) <= 220;
					block_dimensions(3)(1) <= 240;  block_dimensions(19)(1) <= 240;
					block_dimensions(3)(2) <= 280;  block_dimensions(19)(2) <= 240;
					block_dimensions(3)(3) <= 280;  block_dimensions(19)(3) <= 280;
					block_dimensions(4)(0) <= 260;  block_dimensions(20)(0) <= 220;
					block_dimensions(4)(1) <= 320;  block_dimensions(20)(1) <= 320;
					block_dimensions(4)(2) <= 280;  block_dimensions(20)(2) <= 240;
					block_dimensions(4)(3) <= 360;  block_dimensions(20)(3) <= 360;
					block_dimensions(5)(0) <= 260;  block_dimensions(21)(0) <= 220;
					block_dimensions(5)(1) <= 400;  block_dimensions(21)(1) <= 400;
					block_dimensions(5)(2) <= 280;  block_dimensions(21)(2) <= 240;
					block_dimensions(5)(3) <= 440;  block_dimensions(21)(3) <= 440;
					block_dimensions(6)(0) <= 260;  block_dimensions(22)(0) <= 220;
					block_dimensions(6)(1) <= 480;  block_dimensions(22)(1) <= 480;
					block_dimensions(6)(2) <= 280;  block_dimensions(22)(2) <= 240;
					block_dimensions(6)(3) <= 520;  block_dimensions(22)(3) <= 520;
					block_dimensions(7)(0) <= 260;  block_dimensions(23)(0) <= 220;
					block_dimensions(7)(1) <= 560;  block_dimensions(23)(1) <= 560;
					block_dimensions(7)(2) <= 280;  block_dimensions(23)(2) <= 240;
					block_dimensions(7)(3) <= 600;  block_dimensions(23)(3) <= 600;
					block_dimensions(8)(0) <= 240;  block_dimensions(24)(0) <= 200;
					block_dimensions(8)(1) <= 40;   block_dimensions(24)(1) <= 40; 
					block_dimensions(8)(2) <= 260;  block_dimensions(24)(2) <= 220;
					block_dimensions(8)(3) <= 80;   block_dimensions(24)(3) <= 80; 
					block_dimensions(9)(0) <= 240;  block_dimensions(25)(0) <= 200;
					block_dimensions(9)(1) <= 120;  block_dimensions(25)(1) <= 120;
					block_dimensions(9)(2) <= 260;  block_dimensions(25)(2) <= 220;
					block_dimensions(9)(3) <= 160;  block_dimensions(25)(3) <= 160;
					block_dimensions(10)(0) <= 240; block_dimensions(26)(0) <= 200;
                    block_dimensions(10)(1) <= 200; block_dimensions(26)(1) <= 200;                                            
                    block_dimensions(10)(2) <= 260; block_dimensions(26)(2) <= 220;                                            
                    block_dimensions(10)(3) <= 240; block_dimensions(26)(3) <= 240;                                            
                    block_dimensions(11)(0) <= 240; block_dimensions(27)(0) <= 200;                                            
                    block_dimensions(11)(1) <= 280; block_dimensions(27)(1) <= 280;                                            
                    block_dimensions(11)(2) <= 260; block_dimensions(27)(2) <= 220;                                            
                    block_dimensions(11)(3) <= 320; block_dimensions(27)(3) <= 320;                                            
                    block_dimensions(12)(0) <= 240; block_dimensions(28)(0) <= 200;                                            
                    block_dimensions(12)(1) <= 360; block_dimensions(28)(1) <= 360;                                            
                    block_dimensions(12)(2) <= 260; block_dimensions(28)(2) <= 220;                                            
                    block_dimensions(12)(3) <= 400; block_dimensions(28)(3) <= 400;                                            
                    block_dimensions(13)(0) <= 240; block_dimensions(29)(0) <= 200;                                            
                    block_dimensions(13)(1) <= 440; block_dimensions(29)(1) <= 440;                                            
                    block_dimensions(13)(2) <= 260; block_dimensions(29)(2) <= 220;                                            
                    block_dimensions(13)(3) <= 480; block_dimensions(29)(3) <= 480;                                            
                    block_dimensions(14)(0) <= 240; block_dimensions(30)(0) <= 200;                                            
                    block_dimensions(14)(1) <= 520; block_dimensions(30)(1) <= 520;                                            
                    block_dimensions(14)(2) <= 260; block_dimensions(30)(2) <= 220;                                            
                    block_dimensions(14)(3) <= 560; block_dimensions(30)(3) <= 560;                                            
                    block_dimensions(15)(0) <= 240; block_dimensions(31)(0) <= 200;                                            
                    block_dimensions(15)(1) <= 600; block_dimensions(31)(1) <= 600;                                            
                    block_dimensions(15)(2) <= 260; block_dimensions(31)(2) <= 220;                                            
                    block_dimensions(15)(3) <= 640; block_dimensions(31)(3) <= 640;                                            
                                  

                    when "11" =>
					block_dimensions(0)(0) <= 320;  block_dimensions(16)(0) <= 160;
					block_dimensions(0)(1) <= 0;    block_dimensions(16)(1) <= 320;
					block_dimensions(0)(2) <= 360;  block_dimensions(16)(2) <= 200;
					block_dimensions(0)(3) <= 20;   block_dimensions(16)(3) <= 340;
					block_dimensions(1)(0) <= 280;  block_dimensions(17)(0) <= 200;
					block_dimensions(1)(1) <= 20;   block_dimensions(17)(1) <= 340;
					block_dimensions(1)(2) <= 320;  block_dimensions(17)(2) <= 240;
					block_dimensions(1)(3) <= 40;   block_dimensions(17)(3) <= 360;
					block_dimensions(2)(0) <= 240;  block_dimensions(18)(0) <= 240;
					block_dimensions(2)(1) <= 40;   block_dimensions(18)(1) <= 360;
					block_dimensions(2)(2) <= 280;  block_dimensions(18)(2) <= 280;
					block_dimensions(2)(3) <= 60;   block_dimensions(18)(3) <= 380;
					block_dimensions(3)(0) <= 200;  block_dimensions(19)(0) <= 280;
					block_dimensions(3)(1) <= 60;   block_dimensions(19)(1) <= 380;
					block_dimensions(3)(2) <= 240;  block_dimensions(19)(2) <= 320;
					block_dimensions(3)(3) <= 80;   block_dimensions(19)(3) <= 400;
					block_dimensions(4)(0) <= 160;  block_dimensions(20)(0) <= 320;
					block_dimensions(4)(1) <= 80;   block_dimensions(20)(1) <= 400;
					block_dimensions(4)(2) <= 200;  block_dimensions(20)(2) <= 360;
					block_dimensions(4)(3) <= 100;  block_dimensions(20)(3) <= 420;
					block_dimensions(5)(0) <= 120;  block_dimensions(21)(0) <= 280;
					block_dimensions(5)(1) <= 100;  block_dimensions(21)(1) <= 420;
					block_dimensions(5)(2) <= 160;  block_dimensions(21)(2) <= 320;
					block_dimensions(5)(3) <= 120;  block_dimensions(21)(3) <= 440;
					block_dimensions(6)(0) <= 160;  block_dimensions(22)(0) <= 240;
					block_dimensions(6)(1) <= 120;  block_dimensions(22)(1) <= 440;
					block_dimensions(6)(2) <= 200;  block_dimensions(22)(2) <= 280;
					block_dimensions(6)(3) <= 140;  block_dimensions(22)(3) <= 460;
					block_dimensions(7)(0) <= 200;  block_dimensions(23)(0) <= 200;
					block_dimensions(7)(1) <= 140;  block_dimensions(23)(1) <= 460;
					block_dimensions(7)(2) <= 240;  block_dimensions(23)(2) <= 240;
					block_dimensions(7)(3) <= 160;  block_dimensions(23)(3) <= 480;
					block_dimensions(8)(0) <= 240;  block_dimensions(24)(0) <= 160;
					block_dimensions(8)(1) <= 160;  block_dimensions(24)(1) <= 480;
					block_dimensions(8)(2) <= 280;  block_dimensions(24)(2) <= 200;
					block_dimensions(8)(3) <= 180;  block_dimensions(24)(3) <= 500;
					block_dimensions(9)(0) <= 280;  block_dimensions(25)(0) <= 120;
					block_dimensions(9)(1) <= 180;  block_dimensions(25)(1) <= 500;
					block_dimensions(9)(2) <= 320;  block_dimensions(25)(2) <= 160;
					block_dimensions(9)(3) <= 200;  block_dimensions(25)(3) <= 520;
					block_dimensions(10)(0) <= 320; block_dimensions(26)(0) <= 160;
                    block_dimensions(10)(1) <= 200; block_dimensions(26)(1) <= 520;                                            
                    block_dimensions(10)(2) <= 360; block_dimensions(26)(2) <= 200;                                            
                    block_dimensions(10)(3) <= 220; block_dimensions(26)(3) <= 540;                                            
                    block_dimensions(11)(0) <= 280; block_dimensions(27)(0) <= 200;                                            
                    block_dimensions(11)(1) <= 220; block_dimensions(27)(1) <= 540;                                            
                    block_dimensions(11)(2) <= 320; block_dimensions(27)(2) <= 240;                                            
                    block_dimensions(11)(3) <= 240; block_dimensions(27)(3) <= 560;                                            
                    block_dimensions(12)(0) <= 240; block_dimensions(28)(0) <= 240;                                            
                    block_dimensions(12)(1) <= 240; block_dimensions(28)(1) <= 560;                                            
                    block_dimensions(12)(2) <= 280; block_dimensions(28)(2) <= 280;                                            
                    block_dimensions(12)(3) <= 260; block_dimensions(28)(3) <= 580;                                            
                    block_dimensions(13)(0) <= 200; block_dimensions(29)(0) <= 280;                                            
                    block_dimensions(13)(1) <= 260; block_dimensions(29)(1) <= 580;                                            
                    block_dimensions(13)(2) <= 240; block_dimensions(29)(2) <= 320;                                            
                    block_dimensions(13)(3) <= 280; block_dimensions(29)(3) <= 600;                                            
                    block_dimensions(14)(0) <= 160; block_dimensions(30)(0) <= 320;                                            
                    block_dimensions(14)(1) <= 280; block_dimensions(30)(1) <= 600;                                            
                    block_dimensions(14)(2) <= 200; block_dimensions(30)(2) <= 360;                                            
                    block_dimensions(14)(3) <= 300; block_dimensions(30)(3) <= 620;                                            
                    block_dimensions(15)(0) <= 120; block_dimensions(31)(0) <= 280;                                            
                    block_dimensions(15)(1) <= 300; block_dimensions(31)(1) <= 620;                                            
                    block_dimensions(15)(2) <= 160; block_dimensions(31)(2) <= 320;                                            
                    block_dimensions(15)(3) <= 320; block_dimensions(31)(3) <= 640;                                            
                                   
			end case;
		end if;
	end process;
end Behavioral;   